.param d_time = 0.0000000000n