.include "./bisection-params.cir"

.GLOBAL vdd

.param reset_time 	= 1n
.param clk_time 	= 5n

* Supply voltage:
vdd vdd 0 vdd_voltage

* DUT:
.include "./dut.cir"

* Latch inputs:
vp1 reset 	0 pulse (1 0 reset_time 0 0 1 1)
vp2 clk 	0 pulse (0 1 clk_time 	0 0 1 1)
vp3 D  		0 pulse (1 0 d_time		0 0 1 1)
vdc DN 		0 0

* .ic v(x1.a) = 0.5
* .ic v(x1.an) = 0.5

.END
