.include "./bisection-params.cir"

.GLOBAL vdd

* Supply voltage:
vdd vdd 0 vdd_voltage

* DUT:
.include "./dut.cir"

* Latch inputs:
cp1 reset 	0 1
cv2 clk 	0 1
cp3 D  		0 1
cdc DN 		0 1

.include "./ic.cir"

.END
