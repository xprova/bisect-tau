.param d_time = 10.0000000000n