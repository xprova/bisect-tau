.param d_time = 5.0120030872n