.param d_time = 7.5000000000n