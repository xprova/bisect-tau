* Testbench Restart

.GLOBAL vdd

.param reset_time 	= 1n
.param clk_time 	= 5n

* Supply voltage:
vdd vdd 0 vdd_voltage

* DUT:
.include "./dut.cir"

* Latch inputs:
cp1 reset 	0 1
cp2 clk 	0 1
cp3 D  		0 1

.include "./ic.cir"

.END
